library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ram_1_0 is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(6 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_1_0;

architecture Behavioral of ram_1_0 is
   type ram_type is array (0 to 109) of std_logic_vector(15 downto 0);
    signal ram : ram_type := ( 
"1000010101110011", "0000001101101111", "1000010011101111", "1000000001011111", "0000000001101011", "1000011110011111", "1000001011011010", "0000000000000111", "1000001110111000", "1000000101101110", "0000000001101100", "1000001111111110", "0000010001001000", "0000000010001010", "1000010000101010", "1000001010001000", "1000010101000001", "1000011010011001", "0000000001010110", "1000000111000010", "0000000001011101", "1000001001110100", "1000001100010111", "1000000100010100", "1000010111101000","1000010000000101", "1000000001011111", "0000001010110010", "0000000000100110", "1000000010100110", "1000000101000001", "1000001110010000", "1000001111100000", "1000001100110000", "0000000000111010", "1000000000100010", "1000001100011011", "1000001111111011", "0000001000000001", "0000000010101101", "1000001101010010", "1000011101101001", "0000000101010001", "1000000101111101", "1000001000011000", "1000000011111011", "0000001011111111", "0000000100101101", "1000010010011100", "1000000110011001", "1000000101111110", "1000000000101101", "1000001101001100", "1000000001011111", "1000000110011001", "0000000110001000", "1000001110000001", "1000001110001100", "1000011000011111", "0000000110100000", "0000000111111111", "1000000110010011", "0000001001100111", "1000001111000110", "1000000001011010", "1000010101110010", "1000001101010100", "0000000010101100", "1000010101100001", "1000000010111110", "1000001000000010", "0000001001000100", "1000000101110001", "1000011001110111", "1000010001000111", "0000000011100110", "0000001011100010", "1000010000000000", "1000000100101010", "1000001101010000", "0000000011010111", "1000001001011011", "1000001100101110", "1000000000111100", "0000000011000000", "0000000010011111", "1000011101101110", "1000000001110110", "1000000110000011", "1000010111101000", "1000011110010011", "1000000101110011", "1000000001100111", "1000000000100000", "1000000001010001", "1000000100000001", "1000000001101010", "1000000001110111", "0000000111110011", "1000010110100100","1000000101010101", "1000000100100011", "1000000100001001", "1000000110101010", "1000000111011000", "1000000011110000", "1000001010000100", "1000000100010011", "1000001000001110", "1000001011001111");

begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
RAM(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= RAM(conv_integer(a));

end Behavioral;

