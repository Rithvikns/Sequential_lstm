library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_tanh is
    Port ( clk : in std_logic;
we : in std_logic;
a : in STD_LOGIC_vector(15 downto 0);
di : in std_logic_vector(15 downto 0);
do : out std_logic_vector(15 downto 0)
);
end ram_tanh;

architecture Behavioral of ram_tanh is
type mem_array is array (0 to 65535) of std_logic_vector (15 downto 0); 
signal tanh : mem_array := (
0 to 1 => "0000000000000000",
2 to 2 => "0000000000000001",
3 to 3 => "0000000000000010",
4 to 4 => "0000000000000011",
5 to 5 => "0000000000000100",
6 to 6 => "0000000000000101",
7 to 7 => "0000000000000110",
8 to 8 => "0000000000000111",
9 to 9 => "0000000000001000",
10 to 10 => "0000000000001001",
11 to 11 => "0000000000001010",
12 to 12 => "0000000000001011",
13 to 13 => "0000000000001100",
14 to 14 => "0000000000001101",
15 to 15 => "0000000000001110",
16 to 16 => "0000000000001111",
17 to 17 => "0000000000010000",
18 to 18 => "0000000000010001",
19 to 19 => "0000000000010010",
20 to 20 => "0000000000010011",
21 to 21 => "0000000000010100",
22 to 22 => "0000000000010101",
23 to 23 => "0000000000010110",
24 to 24 => "0000000000010111",
25 to 25 => "0000000000011000",
26 to 26 => "0000000000011001",
27 to 27 => "0000000000011010",
28 to 28 => "0000000000011011",
29 to 29 => "0000000000011100",
30 to 30 => "0000000000011101",
31 to 31 => "0000000000011110",
32 to 32 => "0000000000011111",
33 to 33 => "0000000000100000",
34 to 34 => "0000000000100001",
35 to 35 => "0000000000100010",
36 to 36 => "0000000000100011",
37 to 37 => "0000000000100100",
38 to 38 => "0000000000100101",
39 to 39 => "0000000000100110",
40 to 40 => "0000000000100111",
41 to 41 => "0000000000101000",
42 to 42 => "0000000000101001",
43 to 43 => "0000000000101010",
44 to 44 => "0000000000101011",
45 to 45 => "0000000000101100",
46 to 46 => "0000000000101101",
47 to 47 => "0000000000101110",
48 to 48 => "0000000000101111",
49 to 49 => "0000000000110000",
50 to 50 => "0000000000110001",
51 to 51 => "0000000000110010",
52 to 52 => "0000000000110011",
53 to 53 => "0000000000110100",
54 to 54 => "0000000000110101",
55 to 55 => "0000000000110110",
56 to 56 => "0000000000110111",
57 to 57 => "0000000000111000",
58 to 59 => "0000000000111001",
60 to 60 => "0000000000111010",
61 to 61 => "0000000000111011",
62 to 62 => "0000000000111100",
63 to 63 => "0000000000111101",
64 to 64 => "0000000000111110",
65 to 65 => "0000000000111111",
66 to 66 => "0000000001000000",
67 to 67 => "0000000001000001",
68 to 68 => "0000000001000010",
69 to 69 => "0000000001000011",
70 to 70 => "0000000001000100",
71 to 71 => "0000000001000101",
72 to 72 => "0000000001000110",
73 to 73 => "0000000001000111",
74 to 75 => "0000000001001000",
76 to 76 => "0000000001001001",
77 to 77 => "0000000001001010",
78 to 78 => "0000000001001011",
79 to 79 => "0000000001001100",
80 to 80 => "0000000001001101",
81 to 81 => "0000000001001110",
82 to 82 => "0000000001001111",
83 to 83 => "0000000001010000",
84 to 84 => "0000000001010001",
85 to 86 => "0000000001010010",
87 to 87 => "0000000001010011",
88 to 88 => "0000000001010100",
89 to 89 => "0000000001010101",
90 to 90 => "0000000001010110",
91 to 91 => "0000000001010111",
92 to 92 => "0000000001011000",
93 to 94 => "0000000001011001",
95 to 95 => "0000000001011010",
96 to 96 => "0000000001011011",
97 to 97 => "0000000001011100",
98 to 98 => "0000000001011101",
99 to 99 => "0000000001011110",
100 to 100 => "0000000001011111",
101 to 102 => "0000000001100000",
103 to 103 => "0000000001100001",
104 to 104 => "0000000001100010",
105 to 105 => "0000000001100011",
106 to 106 => "0000000001100100",
107 to 107 => "0000000001100101",
108 to 109 => "0000000001100110",
110 to 110 => "0000000001100111",
111 to 111 => "0000000001101000",
112 to 112 => "0000000001101001",
113 to 113 => "0000000001101010",
114 to 115 => "0000000001101011",
116 to 116 => "0000000001101100",
117 to 117 => "0000000001101101",
118 to 118 => "0000000001101110",
119 to 120 => "0000000001101111",
121 to 121 => "0000000001110000",
122 to 122 => "0000000001110001",
123 to 123 => "0000000001110010",
124 to 125 => "0000000001110011",
126 to 126 => "0000000001110100",
127 to 127 => "0000000001110101",
128 to 128 => "0000000001110110",
129 to 130 => "0000000001110111",
131 to 131 => "0000000001111000",
132 to 132 => "0000000001111001",
133 to 134 => "0000000001111010",
135 to 135 => "0000000001111011",
136 to 136 => "0000000001111100",
137 to 137 => "0000000001111101",
138 to 139 => "0000000001111110",
140 to 140 => "0000000001111111",
141 to 141 => "0000000010000000",
142 to 143 => "0000000010000001",
144 to 144 => "0000000010000010",
145 to 146 => "0000000010000011",
147 to 147 => "0000000010000100",
148 to 148 => "0000000010000101",
149 to 150 => "0000000010000110",
151 to 151 => "0000000010000111",
152 to 152 => "0000000010001000",
153 to 154 => "0000000010001001",
155 to 155 => "0000000010001010",
156 to 157 => "0000000010001011",
158 to 158 => "0000000010001100",
159 to 160 => "0000000010001101",
161 to 161 => "0000000010001110",
162 to 162 => "0000000010001111",
163 to 164 => "0000000010010000",
165 to 165 => "0000000010010001",
166 to 167 => "0000000010010010",
168 to 168 => "0000000010010011",
169 to 170 => "0000000010010100",
171 to 171 => "0000000010010101",
172 to 173 => "0000000010010110",
174 to 174 => "0000000010010111",
175 to 176 => "0000000010011000",
177 to 178 => "0000000010011001",
179 to 179 => "0000000010011010",
180 to 181 => "0000000010011011",
182 to 182 => "0000000010011100",
183 to 184 => "0000000010011101",
185 to 186 => "0000000010011110",
187 to 187 => "0000000010011111",
188 to 189 => "0000000010100000",
190 to 190 => "0000000010100001",
191 to 192 => "0000000010100010",
193 to 194 => "0000000010100011",
195 to 196 => "0000000010100100",
197 to 197 => "0000000010100101",
198 to 199 => "0000000010100110",
200 to 201 => "0000000010100111",
202 to 203 => "0000000010101000",
204 to 204 => "0000000010101001",
205 to 206 => "0000000010101010",
207 to 208 => "0000000010101011",
209 to 210 => "0000000010101100",
211 to 212 => "0000000010101101",
213 to 213 => "0000000010101110",
214 to 215 => "0000000010101111",
216 to 217 => "0000000010110000",
218 to 219 => "0000000010110001",
220 to 221 => "0000000010110010",
222 to 223 => "0000000010110011",
224 to 225 => "0000000010110100",
226 to 227 => "0000000010110101",
228 to 229 => "0000000010110110",
230 to 231 => "0000000010110111",
232 to 233 => "0000000010111000",
234 to 235 => "0000000010111001",
236 to 238 => "0000000010111010",
239 to 240 => "0000000010111011",
241 to 242 => "0000000010111100",
243 to 244 => "0000000010111101",
245 to 246 => "0000000010111110",
247 to 249 => "0000000010111111",
250 to 251 => "0000000011000000",
252 to 253 => "0000000011000001",
254 to 256 => "0000000011000010",
257 to 258 => "0000000011000011",
259 to 260 => "0000000011000100",
261 to 263 => "0000000011000101",
264 to 265 => "0000000011000110",
266 to 268 => "0000000011000111",
269 to 271 => "0000000011001000",
272 to 273 => "0000000011001001",
274 to 276 => "0000000011001010",
277 to 279 => "0000000011001011",
280 to 281 => "0000000011001100",
282 to 284 => "0000000011001101",
285 to 287 => "0000000011001110",
288 to 290 => "0000000011001111",
291 to 293 => "0000000011010000",
294 to 296 => "0000000011010001",
297 to 299 => "0000000011010010",
300 to 302 => "0000000011010011",
303 to 305 => "0000000011010100",
306 to 309 => "0000000011010101",
310 to 312 => "0000000011010110",
313 to 315 => "0000000011010111",
316 to 319 => "0000000011011000",
320 to 323 => "0000000011011001",
324 to 326 => "0000000011011010",
327 to 330 => "0000000011011011",
331 to 334 => "0000000011011100",
335 to 338 => "0000000011011101",
339 to 342 => "0000000011011110",
343 to 346 => "0000000011011111",
347 to 350 => "0000000011100000",
351 to 355 => "0000000011100001",
356 to 360 => "0000000011100010",
361 to 364 => "0000000011100011",
365 to 369 => "0000000011100100",
370 to 374 => "0000000011100101",
375 to 380 => "0000000011100110",
381 to 385 => "0000000011100111",
386 to 391 => "0000000011101000",
392 to 397 => "0000000011101001",
398 to 403 => "0000000011101010",
404 to 409 => "0000000011101011",
410 to 416 => "0000000011101100",
417 to 423 => "0000000011101101",
424 to 431 => "0000000011101110",
432 to 439 => "0000000011101111",
440 to 448 => "0000000011110000",
449 to 457 => "0000000011110001",
458 to 466 => "0000000011110010",
467 to 477 => "0000000011110011",
478 to 488 => "0000000011110100",
489 to 501 => "0000000011110101",
502 to 514 => "0000000011110110",
515 to 530 => "0000000011110111",
531 to 547 => "0000000011111000",
548 to 567 => "0000000011111001",
568 to 591 => "0000000011111010",
592 to 620 => "0000000011111011",
621 to 657 => "0000000011111100",
658 to 709 => "0000000011111101",
710 to 798 => "0000000011111110",
799 to 4861 => "0000000011111111",
4862 to 32767 => "0000000100000000",
32768 to 32768 => "0000000000000000",
32769 to 32769 => "1000000000000000",
32770 to 32770 => "1000000000000001",
32771 to 32771 => "1000000000000010",
32772 to 32772 => "1000000000000011",
32773 to 32773 => "1000000000000100",
32774 to 32774 => "1000000000000101",
32775 to 32775 => "1000000000000110",
32776 to 32776 => "1000000000000111",
32777 to 32777 => "1000000000001000",
32778 to 32778 => "1000000000001001",
32779 to 32779 => "1000000000001010",
32780 to 32780 => "1000000000001011",
32781 to 32781 => "1000000000001100",
32782 to 32782 => "1000000000001101",
32783 to 32783 => "1000000000001110",
32784 to 32784 => "1000000000001111",
32785 to 32785 => "1000000000010000",
32786 to 32786 => "1000000000010001",
32787 to 32787 => "1000000000010010",
32788 to 32788 => "1000000000010011",
32789 to 32789 => "1000000000010100",
32790 to 32790 => "1000000000010101",
32791 to 32791 => "1000000000010110",
32792 to 32792 => "1000000000010111",
32793 to 32793 => "1000000000011000",
32794 to 32794 => "1000000000011001",
32795 to 32795 => "1000000000011010",
32796 to 32796 => "1000000000011011",
32797 to 32797 => "1000000000011100",
32798 to 32798 => "1000000000011101",
32799 to 32799 => "1000000000011110",
32800 to 32800 => "1000000000011111",
32801 to 32801 => "1000000000100000",
32802 to 32802 => "1000000000100001",
32803 to 32803 => "1000000000100010",
32804 to 32804 => "1000000000100011",
32805 to 32805 => "1000000000100100",
32806 to 32806 => "1000000000100101",
32807 to 32807 => "1000000000100110",
32808 to 32808 => "1000000000100111",
32809 to 32809 => "1000000000101000",
32810 to 32810 => "1000000000101001",
32811 to 32811 => "1000000000101010",
32812 to 32812 => "1000000000101011",
32813 to 32813 => "1000000000101100",
32814 to 32814 => "1000000000101101",
32815 to 32815 => "1000000000101110",
32816 to 32816 => "1000000000101111",
32817 to 32817 => "1000000000110000",
32818 to 32818 => "1000000000110001",
32819 to 32819 => "1000000000110010",
32820 to 32820 => "1000000000110011",
32821 to 32821 => "1000000000110100",
32822 to 32822 => "1000000000110101",
32823 to 32823 => "1000000000110110",
32824 to 32824 => "1000000000110111",
32825 to 32825 => "1000000000111000",
32826 to 32827 => "1000000000111001",
32828 to 32828 => "1000000000111010",
32829 to 32829 => "1000000000111011",
32830 to 32830 => "1000000000111100",
32831 to 32831 => "1000000000111101",
32832 to 32832 => "1000000000111110",
32833 to 32833 => "1000000000111111",
32834 to 32834 => "1000000001000000",
32835 to 32835 => "1000000001000001",
32836 to 32836 => "1000000001000010",
32837 to 32837 => "1000000001000011",
32838 to 32838 => "1000000001000100",
32839 to 32839 => "1000000001000101",
32840 to 32840 => "1000000001000110",
32841 to 32841 => "1000000001000111",
32842 to 32843 => "1000000001001000",
32844 to 32844 => "1000000001001001",
32845 to 32845 => "1000000001001010",
32846 to 32846 => "1000000001001011",
32847 to 32847 => "1000000001001100",
32848 to 32848 => "1000000001001101",
32849 to 32849 => "1000000001001110",
32850 to 32850 => "1000000001001111",
32851 to 32851 => "1000000001010000",
32852 to 32852 => "1000000001010001",
32853 to 32854 => "1000000001010010",
32855 to 32855 => "1000000001010011",
32856 to 32856 => "1000000001010100",
32857 to 32857 => "1000000001010101",
32858 to 32858 => "1000000001010110",
32859 to 32859 => "1000000001010111",
32860 to 32860 => "1000000001011000",
32861 to 32862 => "1000000001011001",
32863 to 32863 => "1000000001011010",
32864 to 32864 => "1000000001011011",
32865 to 32865 => "1000000001011100",
32866 to 32866 => "1000000001011101",
32867 to 32867 => "1000000001011110",
32868 to 32868 => "1000000001011111",
32869 to 32870 => "1000000001100000",
32871 to 32871 => "1000000001100001",
32872 to 32872 => "1000000001100010",
32873 to 32873 => "1000000001100011",
32874 to 32874 => "1000000001100100",
32875 to 32875 => "1000000001100101",
32876 to 32877 => "1000000001100110",
32878 to 32878 => "1000000001100111",
32879 to 32879 => "1000000001101000",
32880 to 32880 => "1000000001101001",
32881 to 32881 => "1000000001101010",
32882 to 32883 => "1000000001101011",
32884 to 32884 => "1000000001101100",
32885 to 32885 => "1000000001101101",
32886 to 32886 => "1000000001101110",
32887 to 32888 => "1000000001101111",
32889 to 32889 => "1000000001110000",
32890 to 32890 => "1000000001110001",
32891 to 32891 => "1000000001110010",
32892 to 32893 => "1000000001110011",
32894 to 32894 => "1000000001110100",
32895 to 32895 => "1000000001110101",
32896 to 32896 => "1000000001110110",
32897 to 32898 => "1000000001110111",
32899 to 32899 => "1000000001111000",
32900 to 32900 => "1000000001111001",
32901 to 32902 => "1000000001111010",
32903 to 32903 => "1000000001111011",
32904 to 32904 => "1000000001111100",
32905 to 32905 => "1000000001111101",
32906 to 32907 => "1000000001111110",
32908 to 32908 => "1000000001111111",
32909 to 32909 => "1000000010000000",
32910 to 32911 => "1000000010000001",
32912 to 32912 => "1000000010000010",
32913 to 32914 => "1000000010000011",
32915 to 32915 => "1000000010000100",
32916 to 32916 => "1000000010000101",
32917 to 32918 => "1000000010000110",
32919 to 32919 => "1000000010000111",
32920 to 32920 => "1000000010001000",
32921 to 32922 => "1000000010001001",
32923 to 32923 => "1000000010001010",
32924 to 32925 => "1000000010001011",
32926 to 32926 => "1000000010001100",
32927 to 32928 => "1000000010001101",
32929 to 32929 => "1000000010001110",
32930 to 32930 => "1000000010001111",
32931 to 32932 => "1000000010010000",
32933 to 32933 => "1000000010010001",
32934 to 32935 => "1000000010010010",
32936 to 32936 => "1000000010010011",
32937 to 32938 => "1000000010010100",
32939 to 32939 => "1000000010010101",
32940 to 32941 => "1000000010010110",
32942 to 32942 => "1000000010010111",
32943 to 32944 => "1000000010011000",
32945 to 32946 => "1000000010011001",
32947 to 32947 => "1000000010011010",
32948 to 32949 => "1000000010011011",
32950 to 32950 => "1000000010011100",
32951 to 32952 => "1000000010011101",
32953 to 32954 => "1000000010011110",
32955 to 32955 => "1000000010011111",
32956 to 32957 => "1000000010100000",
32958 to 32958 => "1000000010100001",
32959 to 32960 => "1000000010100010",
32961 to 32962 => "1000000010100011",
32963 to 32964 => "1000000010100100",
32965 to 32965 => "1000000010100101",
32966 to 32967 => "1000000010100110",
32968 to 32969 => "1000000010100111",
32970 to 32971 => "1000000010101000",
32972 to 32972 => "1000000010101001",
32973 to 32974 => "1000000010101010",
32975 to 32976 => "1000000010101011",
32977 to 32978 => "1000000010101100",
32979 to 32980 => "1000000010101101",
32981 to 32981 => "1000000010101110",
32982 to 32983 => "1000000010101111",
32984 to 32985 => "1000000010110000",
32986 to 32987 => "1000000010110001",
32988 to 32989 => "1000000010110010",
32990 to 32991 => "1000000010110011",
32992 to 32993 => "1000000010110100",
32994 to 32995 => "1000000010110101",
32996 to 32997 => "1000000010110110",
32998 to 32999 => "1000000010110111",
33000 to 33001 => "1000000010111000",
33002 to 33003 => "1000000010111001",
33004 to 33006 => "1000000010111010",
33007 to 33008 => "1000000010111011",
33009 to 33010 => "1000000010111100",
33011 to 33012 => "1000000010111101",
33013 to 33014 => "1000000010111110",
33015 to 33017 => "1000000010111111",
33018 to 33019 => "1000000011000000",
33020 to 33021 => "1000000011000001",
33022 to 33024 => "1000000011000010",
33025 to 33026 => "1000000011000011",
33027 to 33028 => "1000000011000100",
33029 to 33031 => "1000000011000101",
33032 to 33033 => "1000000011000110",
33034 to 33036 => "1000000011000111",
33037 to 33039 => "1000000011001000",
33040 to 33041 => "1000000011001001",
33042 to 33044 => "1000000011001010",
33045 to 33047 => "1000000011001011",
33048 to 33049 => "1000000011001100",
33050 to 33052 => "1000000011001101",
33053 to 33055 => "1000000011001110",
33056 to 33058 => "1000000011001111",
33059 to 33061 => "1000000011010000",
33062 to 33064 => "1000000011010001",
33065 to 33067 => "1000000011010010",
33068 to 33070 => "1000000011010011",
33071 to 33073 => "1000000011010100",
33074 to 33077 => "1000000011010101",
33078 to 33080 => "1000000011010110",
33081 to 33083 => "1000000011010111",
33084 to 33087 => "1000000011011000",
33088 to 33091 => "1000000011011001",
33092 to 33094 => "1000000011011010",
33095 to 33098 => "1000000011011011",
33099 to 33102 => "1000000011011100",
33103 to 33106 => "1000000011011101",
33107 to 33110 => "1000000011011110",
33111 to 33114 => "1000000011011111",
33115 to 33118 => "1000000011100000",
33119 to 33123 => "1000000011100001",
33124 to 33128 => "1000000011100010",
33129 to 33132 => "1000000011100011",
33133 to 33137 => "1000000011100100",
33138 to 33142 => "1000000011100101",
33143 to 33148 => "1000000011100110",
33149 to 33153 => "1000000011100111",
33154 to 33159 => "1000000011101000",
33160 to 33165 => "1000000011101001",
33166 to 33171 => "1000000011101010",
33172 to 33177 => "1000000011101011",
33178 to 33184 => "1000000011101100",
33185 to 33191 => "1000000011101101",
33192 to 33199 => "1000000011101110",
33200 to 33207 => "1000000011101111",
33208 to 33216 => "1000000011110000",
33217 to 33225 => "1000000011110001",
33226 to 33234 => "1000000011110010",
33235 to 33245 => "1000000011110011",
33246 to 33256 => "1000000011110100",
33257 to 33269 => "1000000011110101",
33270 to 33282 => "1000000011110110",
33283 to 33298 => "1000000011110111",
33299 to 33315 => "1000000011111000",
33316 to 33335 => "1000000011111001",
33336 to 33359 => "1000000011111010",
33360 to 33388 => "1000000011111011",
33389 to 33425 => "1000000011111100",
33426 to 33477 => "1000000011111101",
33478 to 33566 => "1000000011111110",
33567 to 37629 => "1000000011111111",
37630 to 65535 => "1000000100000000");
begin
process (clk)
begin
if (clk'event and clk = '1') then
if (we = '1') then
tanh(conv_integer(a)) <= di;
end if;
end if;
end process;
do <= tanh(conv_integer(a));
end Behavioral;